VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO J1Asic
  CLASS BLOCK ;
  FOREIGN J1Asic ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1960.000 ;
  PIN boardClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END boardClk
  PIN boardClkLocked
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 0.000 712.880 4.000 ;
    END
  END boardClkLocked
  PIN extInt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END extInt[0]
  PIN extInt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END extInt[1]
  PIN extInt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1223.040 0.000 1223.600 4.000 ;
    END
  END extInt[2]
  PIN io_oeb_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1515.360 0.000 1515.920 4.000 ;
    END
  END io_oeb_high[0]
  PIN io_oeb_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1649.760 1956.000 1650.320 1960.000 ;
    END
  END io_oeb_high[1]
  PIN io_oeb_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1622.880 1956.000 1623.440 1960.000 ;
    END
  END io_oeb_high[2]
  PIN io_oeb_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1236.480 0.000 1237.040 4.000 ;
    END
  END io_oeb_high[3]
  PIN io_oeb_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 2032.800 1956.000 2033.360 1960.000 ;
    END
  END io_oeb_high[4]
  PIN io_oeb_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 2479.680 1956.000 2480.240 1960.000 ;
    END
  END io_oeb_high[5]
  PIN io_oeb_high[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1159.200 2800.000 1159.760 ;
    END
  END io_oeb_high[6]
  PIN io_oeb_high[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1579.200 0.000 1579.760 4.000 ;
    END
  END io_oeb_high[7]
  PIN io_oeb_low[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1740.480 0.000 1741.040 4.000 ;
    END
  END io_oeb_low[0]
  PIN io_oeb_low[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1569.120 0.000 1569.680 4.000 ;
    END
  END io_oeb_low[1]
  PIN pmodA_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1307.040 0.000 1307.600 4.000 ;
    END
  END pmodA_oeb[0]
  PIN pmodA_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1404.480 0.000 1405.040 4.000 ;
    END
  END pmodA_oeb[1]
  PIN pmodA_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1458.240 0.000 1458.800 4.000 ;
    END
  END pmodA_oeb[2]
  PIN pmodA_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1767.360 2800.000 1767.920 ;
    END
  END pmodA_oeb[3]
  PIN pmodA_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1659.840 0.000 1660.400 4.000 ;
    END
  END pmodA_oeb[4]
  PIN pmodA_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2503.200 1956.000 2503.760 1960.000 ;
    END
  END pmodA_oeb[5]
  PIN pmodA_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1313.760 0.000 1314.320 4.000 ;
    END
  END pmodA_oeb[6]
  PIN pmodA_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2479.680 0.000 2480.240 4.000 ;
    END
  END pmodA_oeb[7]
  PIN pmodA_read[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1374.240 0.000 1374.800 4.000 ;
    END
  END pmodA_read[0]
  PIN pmodA_read[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1380.960 0.000 1381.520 4.000 ;
    END
  END pmodA_read[1]
  PIN pmodA_read[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1350.720 0.000 1351.280 4.000 ;
    END
  END pmodA_read[2]
  PIN pmodA_read[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 0.000 1354.640 4.000 ;
    END
  END pmodA_read[3]
  PIN pmodA_read[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1303.680 0.000 1304.240 4.000 ;
    END
  END pmodA_read[4]
  PIN pmodA_read[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 0.000 1300.880 4.000 ;
    END
  END pmodA_read[5]
  PIN pmodA_read[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1283.520 0.000 1284.080 4.000 ;
    END
  END pmodA_read[6]
  PIN pmodA_read[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1280.160 0.000 1280.720 4.000 ;
    END
  END pmodA_read[7]
  PIN pmodA_write[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1370.880 0.000 1371.440 4.000 ;
    END
  END pmodA_write[0]
  PIN pmodA_write[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1384.320 0.000 1384.880 4.000 ;
    END
  END pmodA_write[1]
  PIN pmodA_write[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1347.360 0.000 1347.920 4.000 ;
    END
  END pmodA_write[2]
  PIN pmodA_write[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1344.000 0.000 1344.560 4.000 ;
    END
  END pmodA_write[3]
  PIN pmodA_write[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1317.120 0.000 1317.680 4.000 ;
    END
  END pmodA_write[4]
  PIN pmodA_write[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1310.400 0.000 1310.960 4.000 ;
    END
  END pmodA_write[5]
  PIN pmodA_write[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1286.880 0.000 1287.440 4.000 ;
    END
  END pmodA_write[6]
  PIN pmodA_write[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1290.240 0.000 1290.800 4.000 ;
    END
  END pmodA_write[7]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 0.000 675.920 4.000 ;
    END
  END reset
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1149.120 0.000 1149.680 4.000 ;
    END
  END rx
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END tck
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END tdi
  PIN tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 0.000 743.120 4.000 ;
    END
  END tdo
  PIN tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 692.160 4.000 692.720 ;
    END
  END tms
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1135.680 0.000 1136.240 4.000 ;
    END
  END tx
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1944.620 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1944.620 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 2793.280 1945.290 ;
      LAYER Metal2 ;
        RECT 9.100 1955.700 1622.580 1956.000 ;
        RECT 1623.740 1955.700 1649.460 1956.000 ;
        RECT 1650.620 1955.700 2032.500 1956.000 ;
        RECT 2033.660 1955.700 2479.380 1956.000 ;
        RECT 2480.540 1955.700 2502.900 1956.000 ;
        RECT 2504.060 1955.700 2791.460 1956.000 ;
        RECT 9.100 4.300 2791.460 1955.700 ;
        RECT 9.100 3.500 671.700 4.300 ;
        RECT 672.860 3.500 675.060 4.300 ;
        RECT 676.220 3.500 678.420 4.300 ;
        RECT 679.580 3.500 681.780 4.300 ;
        RECT 682.940 3.500 712.020 4.300 ;
        RECT 713.180 3.500 742.260 4.300 ;
        RECT 743.420 3.500 1135.380 4.300 ;
        RECT 1136.540 3.500 1148.820 4.300 ;
        RECT 1149.980 3.500 1222.740 4.300 ;
        RECT 1223.900 3.500 1236.180 4.300 ;
        RECT 1237.340 3.500 1279.860 4.300 ;
        RECT 1281.020 3.500 1283.220 4.300 ;
        RECT 1284.380 3.500 1286.580 4.300 ;
        RECT 1287.740 3.500 1289.940 4.300 ;
        RECT 1291.100 3.500 1300.020 4.300 ;
        RECT 1301.180 3.500 1303.380 4.300 ;
        RECT 1304.540 3.500 1306.740 4.300 ;
        RECT 1307.900 3.500 1310.100 4.300 ;
        RECT 1311.260 3.500 1313.460 4.300 ;
        RECT 1314.620 3.500 1316.820 4.300 ;
        RECT 1317.980 3.500 1343.700 4.300 ;
        RECT 1344.860 3.500 1347.060 4.300 ;
        RECT 1348.220 3.500 1350.420 4.300 ;
        RECT 1351.580 3.500 1353.780 4.300 ;
        RECT 1354.940 3.500 1370.580 4.300 ;
        RECT 1371.740 3.500 1373.940 4.300 ;
        RECT 1375.100 3.500 1380.660 4.300 ;
        RECT 1381.820 3.500 1384.020 4.300 ;
        RECT 1385.180 3.500 1404.180 4.300 ;
        RECT 1405.340 3.500 1457.940 4.300 ;
        RECT 1459.100 3.500 1515.060 4.300 ;
        RECT 1516.220 3.500 1568.820 4.300 ;
        RECT 1569.980 3.500 1578.900 4.300 ;
        RECT 1580.060 3.500 1659.540 4.300 ;
        RECT 1660.700 3.500 1740.180 4.300 ;
        RECT 1741.340 3.500 2479.380 4.300 ;
        RECT 2480.540 3.500 2791.460 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1768.220 2796.000 1944.460 ;
        RECT 4.000 1767.060 2795.700 1768.220 ;
        RECT 4.000 1160.060 2796.000 1767.060 ;
        RECT 4.000 1158.900 2795.700 1160.060 ;
        RECT 4.000 693.020 2796.000 1158.900 ;
        RECT 4.300 691.860 2796.000 693.020 ;
        RECT 4.000 15.540 2796.000 691.860 ;
      LAYER Metal4 ;
        RECT 571.900 17.450 636.340 1916.230 ;
        RECT 638.540 17.450 713.140 1916.230 ;
        RECT 715.340 17.450 789.940 1916.230 ;
        RECT 792.140 17.450 866.740 1916.230 ;
        RECT 868.940 17.450 943.540 1916.230 ;
        RECT 945.740 17.450 1020.340 1916.230 ;
        RECT 1022.540 17.450 1097.140 1916.230 ;
        RECT 1099.340 17.450 1173.940 1916.230 ;
        RECT 1176.140 17.450 1250.740 1916.230 ;
        RECT 1252.940 17.450 1327.540 1916.230 ;
        RECT 1329.740 17.450 1404.340 1916.230 ;
        RECT 1406.540 17.450 1481.140 1916.230 ;
        RECT 1483.340 17.450 1557.940 1916.230 ;
        RECT 1560.140 17.450 1634.740 1916.230 ;
        RECT 1636.940 17.450 1711.540 1916.230 ;
        RECT 1713.740 17.450 1788.340 1916.230 ;
        RECT 1790.540 17.450 1865.140 1916.230 ;
        RECT 1867.340 17.450 1941.940 1916.230 ;
        RECT 1944.140 17.450 2018.740 1916.230 ;
        RECT 2020.940 17.450 2095.540 1916.230 ;
        RECT 2097.740 17.450 2172.340 1916.230 ;
        RECT 2174.540 17.450 2249.140 1916.230 ;
        RECT 2251.340 17.450 2325.940 1916.230 ;
        RECT 2328.140 17.450 2402.740 1916.230 ;
        RECT 2404.940 17.450 2479.540 1916.230 ;
        RECT 2481.740 17.450 2499.700 1916.230 ;
  END
END J1Asic
END LIBRARY

