magic
tech gf180mcuD
magscale 1 5
timestamp 1702222513
<< obsm1 >>
rect 672 855 279328 194529
<< metal2 >>
rect 162288 195600 162344 196000
rect 164976 195600 165032 196000
rect 203280 195600 203336 196000
rect 247968 195600 248024 196000
rect 250320 195600 250376 196000
rect 0 0 56 400
rect 336 0 392 400
rect 67200 0 67256 400
rect 67536 0 67592 400
rect 67872 0 67928 400
rect 68208 0 68264 400
rect 71232 0 71288 400
rect 74256 0 74312 400
rect 113568 0 113624 400
rect 114912 0 114968 400
rect 122304 0 122360 400
rect 123648 0 123704 400
rect 128016 0 128072 400
rect 128352 0 128408 400
rect 128688 0 128744 400
rect 129024 0 129080 400
rect 130032 0 130088 400
rect 130368 0 130424 400
rect 130704 0 130760 400
rect 131040 0 131096 400
rect 131376 0 131432 400
rect 131712 0 131768 400
rect 134400 0 134456 400
rect 134736 0 134792 400
rect 135072 0 135128 400
rect 135408 0 135464 400
rect 137088 0 137144 400
rect 137424 0 137480 400
rect 138096 0 138152 400
rect 138432 0 138488 400
rect 140448 0 140504 400
rect 145824 0 145880 400
rect 151536 0 151592 400
rect 156912 0 156968 400
rect 157920 0 157976 400
rect 165984 0 166040 400
rect 174048 0 174104 400
rect 247968 0 248024 400
<< obsm2 >>
rect 910 195570 162258 195600
rect 162374 195570 164946 195600
rect 165062 195570 203250 195600
rect 203366 195570 247938 195600
rect 248054 195570 250290 195600
rect 250406 195570 279146 195600
rect 910 430 279146 195570
rect 910 350 67170 430
rect 67286 350 67506 430
rect 67622 350 67842 430
rect 67958 350 68178 430
rect 68294 350 71202 430
rect 71318 350 74226 430
rect 74342 350 113538 430
rect 113654 350 114882 430
rect 114998 350 122274 430
rect 122390 350 123618 430
rect 123734 350 127986 430
rect 128102 350 128322 430
rect 128438 350 128658 430
rect 128774 350 128994 430
rect 129110 350 130002 430
rect 130118 350 130338 430
rect 130454 350 130674 430
rect 130790 350 131010 430
rect 131126 350 131346 430
rect 131462 350 131682 430
rect 131798 350 134370 430
rect 134486 350 134706 430
rect 134822 350 135042 430
rect 135158 350 135378 430
rect 135494 350 137058 430
rect 137174 350 137394 430
rect 137510 350 138066 430
rect 138182 350 138402 430
rect 138518 350 140418 430
rect 140534 350 145794 430
rect 145910 350 151506 430
rect 151622 350 156882 430
rect 156998 350 157890 430
rect 158006 350 165954 430
rect 166070 350 174018 430
rect 174134 350 247938 430
rect 248054 350 279146 430
<< metal3 >>
rect 279600 176736 280000 176792
rect 279600 115920 280000 115976
rect 0 69216 400 69272
<< obsm3 >>
rect 400 176822 279600 194446
rect 400 176706 279570 176822
rect 400 116006 279600 176706
rect 400 115890 279570 116006
rect 400 69302 279600 115890
rect 430 69186 279600 69302
rect 400 1554 279600 69186
<< metal4 >>
rect 2224 1538 2384 194462
rect 9904 1538 10064 194462
rect 17584 1538 17744 194462
rect 25264 1538 25424 194462
rect 32944 1538 33104 194462
rect 40624 1538 40784 194462
rect 48304 1538 48464 194462
rect 55984 1538 56144 194462
rect 63664 1538 63824 194462
rect 71344 1538 71504 194462
rect 79024 1538 79184 194462
rect 86704 1538 86864 194462
rect 94384 1538 94544 194462
rect 102064 1538 102224 194462
rect 109744 1538 109904 194462
rect 117424 1538 117584 194462
rect 125104 1538 125264 194462
rect 132784 1538 132944 194462
rect 140464 1538 140624 194462
rect 148144 1538 148304 194462
rect 155824 1538 155984 194462
rect 163504 1538 163664 194462
rect 171184 1538 171344 194462
rect 178864 1538 179024 194462
rect 186544 1538 186704 194462
rect 194224 1538 194384 194462
rect 201904 1538 202064 194462
rect 209584 1538 209744 194462
rect 217264 1538 217424 194462
rect 224944 1538 225104 194462
rect 232624 1538 232784 194462
rect 240304 1538 240464 194462
rect 247984 1538 248144 194462
rect 255664 1538 255824 194462
rect 263344 1538 263504 194462
rect 271024 1538 271184 194462
rect 278704 1538 278864 194462
<< obsm4 >>
rect 57190 1745 63634 191623
rect 63854 1745 71314 191623
rect 71534 1745 78994 191623
rect 79214 1745 86674 191623
rect 86894 1745 94354 191623
rect 94574 1745 102034 191623
rect 102254 1745 109714 191623
rect 109934 1745 117394 191623
rect 117614 1745 125074 191623
rect 125294 1745 132754 191623
rect 132974 1745 140434 191623
rect 140654 1745 148114 191623
rect 148334 1745 155794 191623
rect 156014 1745 163474 191623
rect 163694 1745 171154 191623
rect 171374 1745 178834 191623
rect 179054 1745 186514 191623
rect 186734 1745 194194 191623
rect 194414 1745 201874 191623
rect 202094 1745 209554 191623
rect 209774 1745 217234 191623
rect 217454 1745 224914 191623
rect 225134 1745 232594 191623
rect 232814 1745 240274 191623
rect 240494 1745 247954 191623
rect 248174 1745 249970 191623
<< labels >>
rlabel metal2 s 67200 0 67256 400 6 boardClk
port 1 nsew signal input
rlabel metal2 s 71232 0 71288 400 6 boardClkLocked
port 2 nsew signal input
rlabel metal2 s 0 0 56 400 6 extInt[0]
port 3 nsew signal input
rlabel metal2 s 336 0 392 400 6 extInt[1]
port 4 nsew signal input
rlabel metal2 s 122304 0 122360 400 6 extInt[2]
port 5 nsew signal input
rlabel metal2 s 151536 0 151592 400 6 io_oeb_high[0]
port 6 nsew signal output
rlabel metal2 s 164976 195600 165032 196000 6 io_oeb_high[1]
port 7 nsew signal output
rlabel metal2 s 162288 195600 162344 196000 6 io_oeb_high[2]
port 8 nsew signal output
rlabel metal2 s 123648 0 123704 400 6 io_oeb_high[3]
port 9 nsew signal output
rlabel metal2 s 203280 195600 203336 196000 6 io_oeb_high[4]
port 10 nsew signal output
rlabel metal2 s 247968 195600 248024 196000 6 io_oeb_high[5]
port 11 nsew signal output
rlabel metal3 s 279600 115920 280000 115976 6 io_oeb_high[6]
port 12 nsew signal output
rlabel metal2 s 157920 0 157976 400 6 io_oeb_high[7]
port 13 nsew signal output
rlabel metal2 s 174048 0 174104 400 6 io_oeb_low[0]
port 14 nsew signal output
rlabel metal2 s 156912 0 156968 400 6 io_oeb_low[1]
port 15 nsew signal output
rlabel metal2 s 130704 0 130760 400 6 pmodA_oeb[0]
port 16 nsew signal output
rlabel metal2 s 140448 0 140504 400 6 pmodA_oeb[1]
port 17 nsew signal output
rlabel metal2 s 145824 0 145880 400 6 pmodA_oeb[2]
port 18 nsew signal output
rlabel metal3 s 279600 176736 280000 176792 6 pmodA_oeb[3]
port 19 nsew signal output
rlabel metal2 s 165984 0 166040 400 6 pmodA_oeb[4]
port 20 nsew signal output
rlabel metal2 s 250320 195600 250376 196000 6 pmodA_oeb[5]
port 21 nsew signal output
rlabel metal2 s 131376 0 131432 400 6 pmodA_oeb[6]
port 22 nsew signal output
rlabel metal2 s 247968 0 248024 400 6 pmodA_oeb[7]
port 23 nsew signal output
rlabel metal2 s 137424 0 137480 400 6 pmodA_read[0]
port 24 nsew signal input
rlabel metal2 s 138096 0 138152 400 6 pmodA_read[1]
port 25 nsew signal input
rlabel metal2 s 135072 0 135128 400 6 pmodA_read[2]
port 26 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 pmodA_read[3]
port 27 nsew signal input
rlabel metal2 s 130368 0 130424 400 6 pmodA_read[4]
port 28 nsew signal input
rlabel metal2 s 130032 0 130088 400 6 pmodA_read[5]
port 29 nsew signal input
rlabel metal2 s 128352 0 128408 400 6 pmodA_read[6]
port 30 nsew signal input
rlabel metal2 s 128016 0 128072 400 6 pmodA_read[7]
port 31 nsew signal input
rlabel metal2 s 137088 0 137144 400 6 pmodA_write[0]
port 32 nsew signal output
rlabel metal2 s 138432 0 138488 400 6 pmodA_write[1]
port 33 nsew signal output
rlabel metal2 s 134736 0 134792 400 6 pmodA_write[2]
port 34 nsew signal output
rlabel metal2 s 134400 0 134456 400 6 pmodA_write[3]
port 35 nsew signal output
rlabel metal2 s 131712 0 131768 400 6 pmodA_write[4]
port 36 nsew signal output
rlabel metal2 s 131040 0 131096 400 6 pmodA_write[5]
port 37 nsew signal output
rlabel metal2 s 128688 0 128744 400 6 pmodA_write[6]
port 38 nsew signal output
rlabel metal2 s 129024 0 129080 400 6 pmodA_write[7]
port 39 nsew signal output
rlabel metal2 s 67536 0 67592 400 6 reset
port 40 nsew signal input
rlabel metal2 s 114912 0 114968 400 6 rx
port 41 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 tck
port 42 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 tdi
port 43 nsew signal input
rlabel metal2 s 74256 0 74312 400 6 tdo
port 44 nsew signal output
rlabel metal3 s 0 69216 400 69272 6 tms
port 45 nsew signal input
rlabel metal2 s 113568 0 113624 400 6 tx
port 46 nsew signal output
rlabel metal4 s 2224 1538 2384 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 194462 6 vdd
port 47 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 194462 6 vss
port 48 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 194462 6 vss
port 48 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 280000 196000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 71240238
string GDS_FILE /home/moss/eda_tools_gf180_new/caravel_user_project/openlane/J1Asic/runs/23_12_10_14_39/results/signoff/J1Asic.magic.gds
string GDS_START 606712
<< end >>

