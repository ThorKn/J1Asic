VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO J1Asic
  CLASS BLOCK ;
  FOREIGN J1Asic ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1960.000 ;
  PIN boardClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END boardClk
  PIN boardClkLocked
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 0.000 938.000 4.000 ;
    END
  END boardClkLocked
  PIN extInt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END extInt[0]
  PIN extInt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END extInt[1]
  PIN extInt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1559.040 0.000 1559.600 4.000 ;
    END
  END extInt[2]
  PIN io_oeb_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1337.280 0.000 1337.840 4.000 ;
    END
  END io_oeb_high[0]
  PIN io_oeb_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1115.520 0.000 1116.080 4.000 ;
    END
  END io_oeb_high[1]
  PIN io_oeb_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1871.520 1956.000 1872.080 1960.000 ;
    END
  END io_oeb_high[2]
  PIN io_oeb_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1596.000 1956.000 1596.560 1960.000 ;
    END
  END io_oeb_high[3]
  PIN io_oeb_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1357.440 0.000 1358.000 4.000 ;
    END
  END io_oeb_high[4]
  PIN io_oeb_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1737.120 0.000 1737.680 4.000 ;
    END
  END io_oeb_high[5]
  PIN io_oeb_high[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1246.560 0.000 1247.120 4.000 ;
    END
  END io_oeb_high[6]
  PIN io_oeb_high[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 1512.000 0.000 1512.560 4.000 ;
    END
  END io_oeb_high[7]
  PIN io_oeb_low[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 0.000 1663.760 4.000 ;
    END
  END io_oeb_low[0]
  PIN io_oeb_low[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1733.760 1956.000 1734.320 1960.000 ;
    END
  END io_oeb_low[1]
  PIN pmodA_read[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1424.640 0.000 1425.200 4.000 ;
    END
  END pmodA_read[0]
  PIN pmodA_read[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1404.480 0.000 1405.040 4.000 ;
    END
  END pmodA_read[1]
  PIN pmodA_read[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1401.120 0.000 1401.680 4.000 ;
    END
  END pmodA_read[2]
  PIN pmodA_read[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1377.600 0.000 1378.160 4.000 ;
    END
  END pmodA_read[3]
  PIN pmodA_read[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1384.320 0.000 1384.880 4.000 ;
    END
  END pmodA_read[4]
  PIN pmodA_read[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1350.720 0.000 1351.280 4.000 ;
    END
  END pmodA_read[5]
  PIN pmodA_read[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 0.000 1354.640 4.000 ;
    END
  END pmodA_read[6]
  PIN pmodA_read[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1360.800 0.000 1361.360 4.000 ;
    END
  END pmodA_read[7]
  PIN pmodA_writeEnable[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1417.920 0.000 1418.480 4.000 ;
    END
  END pmodA_writeEnable[0]
  PIN pmodA_writeEnable[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1394.400 0.000 1394.960 4.000 ;
    END
  END pmodA_writeEnable[1]
  PIN pmodA_writeEnable[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1391.040 0.000 1391.600 4.000 ;
    END
  END pmodA_writeEnable[2]
  PIN pmodA_writeEnable[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1370.880 0.000 1371.440 4.000 ;
    END
  END pmodA_writeEnable[3]
  PIN pmodA_writeEnable[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1414.560 0.000 1415.120 4.000 ;
    END
  END pmodA_writeEnable[4]
  PIN pmodA_writeEnable[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1387.680 0.000 1388.240 4.000 ;
    END
  END pmodA_writeEnable[5]
  PIN pmodA_writeEnable[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1344.000 0.000 1344.560 4.000 ;
    END
  END pmodA_writeEnable[6]
  PIN pmodA_writeEnable[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1411.200 0.000 1411.760 4.000 ;
    END
  END pmodA_writeEnable[7]
  PIN pmodA_write[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1421.280 0.000 1421.840 4.000 ;
    END
  END pmodA_write[0]
  PIN pmodA_write[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1407.840 0.000 1408.400 4.000 ;
    END
  END pmodA_write[1]
  PIN pmodA_write[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1397.760 0.000 1398.320 4.000 ;
    END
  END pmodA_write[2]
  PIN pmodA_write[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1374.240 0.000 1374.800 4.000 ;
    END
  END pmodA_write[3]
  PIN pmodA_write[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1380.960 0.000 1381.520 4.000 ;
    END
  END pmodA_write[4]
  PIN pmodA_write[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1347.360 0.000 1347.920 4.000 ;
    END
  END pmodA_write[5]
  PIN pmodA_write[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1364.160 0.000 1364.720 4.000 ;
    END
  END pmodA_write[6]
  PIN pmodA_write[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 0.000 1368.080 4.000 ;
    END
  END pmodA_write[7]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 0.000 927.920 4.000 ;
    END
  END reset
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1223.040 0.000 1223.600 4.000 ;
    END
  END rx
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 0.000 753.200 4.000 ;
    END
  END tck
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 0.000 948.080 4.000 ;
    END
  END tdi
  PIN tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1041.600 0.000 1042.160 4.000 ;
    END
  END tdo
  PIN tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 0.000 897.680 4.000 ;
    END
  END tms
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1229.760 0.000 1230.320 4.000 ;
    END
  END tx
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1944.620 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1944.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1944.620 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 2793.280 1944.620 ;
      LAYER Metal2 ;
        RECT 22.380 1955.700 1595.700 1956.000 ;
        RECT 1596.860 1955.700 1733.460 1956.000 ;
        RECT 1734.620 1955.700 1871.220 1956.000 ;
        RECT 1872.380 1955.700 2788.500 1956.000 ;
        RECT 22.380 4.300 2788.500 1955.700 ;
        RECT 22.380 3.500 671.700 4.300 ;
        RECT 672.860 3.500 752.340 4.300 ;
        RECT 753.500 3.500 896.820 4.300 ;
        RECT 897.980 3.500 927.060 4.300 ;
        RECT 928.220 3.500 937.140 4.300 ;
        RECT 938.300 3.500 947.220 4.300 ;
        RECT 948.380 3.500 1041.300 4.300 ;
        RECT 1042.460 3.500 1115.220 4.300 ;
        RECT 1116.380 3.500 1222.740 4.300 ;
        RECT 1223.900 3.500 1229.460 4.300 ;
        RECT 1230.620 3.500 1246.260 4.300 ;
        RECT 1247.420 3.500 1336.980 4.300 ;
        RECT 1338.140 3.500 1343.700 4.300 ;
        RECT 1344.860 3.500 1347.060 4.300 ;
        RECT 1348.220 3.500 1350.420 4.300 ;
        RECT 1351.580 3.500 1353.780 4.300 ;
        RECT 1354.940 3.500 1357.140 4.300 ;
        RECT 1358.300 3.500 1360.500 4.300 ;
        RECT 1361.660 3.500 1363.860 4.300 ;
        RECT 1365.020 3.500 1367.220 4.300 ;
        RECT 1368.380 3.500 1370.580 4.300 ;
        RECT 1371.740 3.500 1373.940 4.300 ;
        RECT 1375.100 3.500 1377.300 4.300 ;
        RECT 1378.460 3.500 1380.660 4.300 ;
        RECT 1381.820 3.500 1384.020 4.300 ;
        RECT 1385.180 3.500 1387.380 4.300 ;
        RECT 1388.540 3.500 1390.740 4.300 ;
        RECT 1391.900 3.500 1394.100 4.300 ;
        RECT 1395.260 3.500 1397.460 4.300 ;
        RECT 1398.620 3.500 1400.820 4.300 ;
        RECT 1401.980 3.500 1404.180 4.300 ;
        RECT 1405.340 3.500 1407.540 4.300 ;
        RECT 1408.700 3.500 1410.900 4.300 ;
        RECT 1412.060 3.500 1414.260 4.300 ;
        RECT 1415.420 3.500 1417.620 4.300 ;
        RECT 1418.780 3.500 1420.980 4.300 ;
        RECT 1422.140 3.500 1424.340 4.300 ;
        RECT 1425.500 3.500 1511.700 4.300 ;
        RECT 1512.860 3.500 1558.740 4.300 ;
        RECT 1559.900 3.500 1662.900 4.300 ;
        RECT 1664.060 3.500 1736.820 4.300 ;
        RECT 1737.980 3.500 2788.500 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 15.540 2788.550 1944.460 ;
      LAYER Metal4 ;
        RECT 454.300 17.450 482.740 1823.830 ;
        RECT 484.940 17.450 559.540 1823.830 ;
        RECT 561.740 17.450 636.340 1823.830 ;
        RECT 638.540 17.450 713.140 1823.830 ;
        RECT 715.340 17.450 789.940 1823.830 ;
        RECT 792.140 17.450 866.740 1823.830 ;
        RECT 868.940 17.450 943.540 1823.830 ;
        RECT 945.740 17.450 1020.340 1823.830 ;
        RECT 1022.540 17.450 1097.140 1823.830 ;
        RECT 1099.340 17.450 1173.940 1823.830 ;
        RECT 1176.140 17.450 1250.740 1823.830 ;
        RECT 1252.940 17.450 1327.540 1823.830 ;
        RECT 1329.740 17.450 1404.340 1823.830 ;
        RECT 1406.540 17.450 1481.140 1823.830 ;
        RECT 1483.340 17.450 1557.940 1823.830 ;
        RECT 1560.140 17.450 1634.740 1823.830 ;
        RECT 1636.940 17.450 1711.540 1823.830 ;
        RECT 1713.740 17.450 1788.340 1823.830 ;
        RECT 1790.540 17.450 1865.140 1823.830 ;
        RECT 1867.340 17.450 1941.940 1823.830 ;
        RECT 1944.140 17.450 2018.740 1823.830 ;
        RECT 2020.940 17.450 2095.540 1823.830 ;
        RECT 2097.740 17.450 2172.340 1823.830 ;
        RECT 2174.540 17.450 2249.140 1823.830 ;
        RECT 2251.340 17.450 2325.940 1823.830 ;
        RECT 2328.140 17.450 2402.740 1823.830 ;
        RECT 2404.940 17.450 2452.100 1823.830 ;
  END
END J1Asic
END LIBRARY

